--------------------------------------------------------------------------------
-- Company: UVigo
-- Engineer: Jacobo Cabaleiro
--
-- Create Date:    
-- Design Name:    
-- Module Name:    cordic - beh
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
-- | *** SPECS ***
-- | Latency: 8 cycles
-- | Throughoutput: 1 sample / 8 cycles
-- |
-- | *** BRIEF DESCRIPTION ***
-- | Cordic based sequential engine for generating sin and cosine values from radian 
-- | angles.
-- |
-- | *** DESCRIPTION ***
-- | Sequential iterative cordic based sin / cos calculator. Works on clock
-- | rising edge and includes a synchronous reset signal so it can be put on a known
-- | state (done state).
-- |
-- | ** Ports **
-- | * Inputs *
-- | -> CLK
-- | -> RST: synchronous reset
-- | -> RUN: run/done iface run signal. See below for description
-- | -> ANGLE: input angle, in radians
-- | * Outputs *
-- | -> SIN: sin value for given input angle
-- | -> COS: cos value for given input angle
-- | -> DONE: run/done iface done signal. See below for description
-- |
-- *** RUN / DONE interface ***
-- // THIS SHOULD BE USED AS THE RUN / DONE MAIN SPECIFICATION //
-- Runs on rising edge of clocks. If run signal is low, cordic stays in a "done" state
-- giving the last calculated sin / cos values. If run is pulled up, next cicle the 
-- engine starts calculating the sin & cos for the angle found in its input.
--
-- Run can the be pulled down again as engine will be calculating till it obtains the value
-- (it takes it 8 cycles). In the CYCLE THE ELEMENT KNOWS WILL HAVE THE VALUE
-- READY, sets the DONE port high again. So, BEFORE the next rising edge, the
-- value is ready and stable in its output. This way (1 "cycle advance" in announcing the result is ready) an
-- | optimal chaining of repetitive calcs can be done without otherwise loosing at least one
-- | clock cycle.
--
-- Todo:
-- * Everything should be parametrized, even the number of output precision
-- bits (which in turn changes latency)
--
-- Dependencies:
-- 
-- Revision:
-- MARK -> revision 0.03 has been tested. Works OK. Small problems with
-- precision appear near 0 radians
-- Revision 0.03 - Counter reset is now synchronous (UNTESTED)
-- Revision 0.02 - New state machine (TESTED)
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use WORK.COMMON.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cordic is
        -- rev 0.03
	generic (
		width : natural := PIPELINE_WIDTH
	);
	port (
		clk, rst, run : in std_logic;
		angle : in std_logic_vector(width - 1 downto 0); -- In RADIANS!
		sin, cos : out std_logic_vector(width - 1 downto 0);
		done : out std_logic
	);
end cordic;

architecture beh of cordic is
	type state_t is (
		ST_DONE, ST_INIT, ST_RUNNING, ST_LAST
	);

	signal st : state_t; -- Se podr�a hacer con una variable compartida, aunque debido al posible comportamiento no determinista se prefiere simular (como en la realidad) mediante una se�al
	signal step : std_logic_vector(2 downto 0);

	-- Control signas (generated by FSM)
	signal init, save : std_logic;

	-- Cordic interconnect signals
	signal x0, y0 : std_logic_vector(width - 1 downto 0);
	signal gt_hPI_s, lt_mhPI_s : std_logic;
	signal z_add_sub_op : std_logic;
	signal x_mux_out, y_mux_out, z_mux_out : std_logic_vector(width - 1 downto 0);
	signal z_delta_mux_out, atan_lut_out : std_logic_vector(width - 1 downto 0);
	signal x_reg_out, y_reg_out, z_reg_out : std_logic_vector(width - 1 downto 0);
	signal x_add_sub_out, y_add_sub_out, z_add_sub_out : std_logic_vector(width - 1 downto 0);
	signal x_shift_out, y_shift_out : std_logic_vector(width - 1 downto 0);

	alias z_msb : std_logic is z_reg_out(width - 1);
	signal n_z_msb : std_logic;

	-- Components
	component add_sub is
		generic (
			width : natural := PIPELINE_WIDTH
		);
		port (
			a, b: in std_logic_vector(width - 1 downto 0);
			add_nsub : in std_logic;
			o: out std_logic_vector(width - 1 downto 0);
			f_ov, f_z: out std_logic
		);
	end component;

	component reg is
		generic (
			width : natural := PIPELINE_WIDTH
		);
		port (
			clk, we, rst : in std_logic;
			i : in std_logic_vector (width - 1 downto 0);
			o : out std_logic_vector (width - 1 downto 0)
		);
	end component;

	component signed_r_shifter is
		generic (
			width : natural := PIPELINE_WIDTH;
			width_dir_bits : natural := PIPELINE_WIDTH_DIR_BITS
		);
		port (
			i : in std_logic_vector(width - 1 downto 0);
			n : in std_logic_vector(width_dir_bits - 1 downto 0);
			o : out std_logic_vector(width - 1 downto 0)
		);
	end component;

	component k_lt_comp is
		generic (
			width : natural := PIPELINE_WIDTH;
			k : pipeline_integer := 0
		);
		port (
			a : in std_logic_vector(width - 1 downto 0);
			a_lt_k : out std_logic
		);
	end component;

	component k_gt_comp is
		generic (
			width : natural := PIPELINE_WIDTH;
			k : pipeline_integer := 0
		);
		port (
			a : in std_logic_vector(width - 1 downto 0);
			a_gt_k : out std_logic
		);
	end component;

	component cordic_elem_init is
		generic (
			width : natural := PIPELINE_WIDTH
		);
		port (
			gt_hPI, lt_mhPI : in std_logic;
			x_init_val, y_init_val : out std_logic_vector(width - 1 downto 0)
		);	
	end component;

	component cord_atan_lut is
		port (
			addr : in std_logic_vector(2 downto 0);
			angle : out std_logic_vector(15 downto 0)
		);
	end component;
begin
	-- Instanciaciones de los componentes
	lt_comp : k_lt_comp
		generic map (
			k => MINUS_HALF_PI_FX316
		)
		port map (
			a => angle,
			a_lt_k => lt_mhPI_s
		);

	gt_comp : k_gt_comp
		generic map (
			k => HALF_PI_FX316
		)
		port map (
			a => angle,
			a_gt_k => gt_hPI_s
		);

	elem_init : cordic_elem_init
		port map (
			gt_hPI => gt_hPI_s,
			lt_mhPI => lt_mhPI_s,
			x_init_val => x0,
			y_init_val => y0
		);

	x_add_sub : add_sub
		port map (
			-- ENTRADAS
			a => x_reg_out,
			b => y_shift_out,
			add_nsub => z_msb,
			-- SALIDAS
			o => x_add_sub_out,
                        -- Unconnected
                        f_ov => open,
                        f_z => open
		);

	y_add_sub : add_sub
		port map (
			-- ENTRADAS
			a => y_reg_out,
			b => x_shift_out,
			add_nsub => n_z_msb,
			-- SALIDAS
			o => y_add_sub_out,
                        -- Unconnected
                        f_ov => open,
                        f_z => open
		);

	z_add_sub : add_sub
		port map (
			-- ENTRADAS
			a => z_mux_out,
			b => z_delta_mux_out,
			add_nsub => z_add_sub_op,
			-- SALIDS
			o => z_add_sub_out
		);

	x_reg : reg
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => x_mux_out,
			-- SALIDAS
			o => x_reg_out
		);

	y_reg : reg
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => y_mux_out,
			-- SALIDAS
			o => y_reg_out
		);

	z_reg : reg
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => z_add_sub_out,
			-- SALIDAS
			o => z_reg_out
		);

	cos_reg : reg
		port map (
			-- ENTRADAS
			clk => clk, we => save, rst => rst,
			i => x_add_sub_out,
			-- SALIDAS
			o => cos
		);

	sin_reg : reg
		port map (
			-- ENTRADAS
			clk => clk, we => save, rst => rst,
			i => y_add_sub_out,
			-- SALIDAS
			o => sin
		);

	x_shifter : signed_r_shifter
		port map (
			-- ENTRADAS
			i => x_reg_out,
			n(3) => '0', n(2 downto 0) => step,
			-- SALIDAS
			o => x_shift_out
		);

	y_shifter : signed_r_shifter
		port map (
			-- ENTRADAS
			i => y_reg_out,
			n(3) => '0', n(2 downto 0) => step,
			-- SALIDAS
			o => y_shift_out
		);

	atan_lut : cord_atan_lut
		port map (
			addr => step,
			angle => atan_lut_out
		);

	state_ctrl : process(clk, run, rst)
	begin
		if (rising_edge(clk)) then
			if (rst = '1') then
				st <= ST_DONE;
			else
				case st is
					when ST_DONE =>
						if (run = '1') then
							st <= ST_INIT;
						else
							st <= ST_DONE;
						end if;
					when ST_INIT =>
						st <= ST_RUNNING;
					when ST_RUNNING =>
						if (step = "110") then
							st <= ST_LAST;
						else
							st <= ST_RUNNING;
						end if;
					when ST_LAST =>
                                                st <= ST_DONE;
					when others =>
						assert true
							report "Unkown state!!! Should not happen!!!"
							severity error;
						st <= st;
				end case;
			end if;
		end if;
	end process state_ctrl;

	step_counter : process(clk)
		subtype step_counter_t is natural range 0 to 7;
		variable step_counter : step_counter_t;
	begin
		if (rising_edge(clk)) then
			if (init = '1') then
				step_counter := 0;
			else
				-- Just fold if I'm out of range
				if (step_counter = step_counter_t'high) then
					step_counter := 0;
				else
					step_counter := step_counter + 1;
				end if;
			end if;
		end if;
		step <= std_logic_vector(to_unsigned(step_counter,3));
	end process;

	signals_gen : process(st)
	begin
		case st is
			when ST_DONE =>
				init <= '0';
				save <= '0';
				done <= '1';
			when ST_INIT =>
				init <= '1';
				save <= '0';
				done <= '0';
			when ST_RUNNING =>
				init <= '0';
				save <= '0';
				done <= '0';
			when ST_LAST =>
				save <= '1';
				init <= '0';
				done <= '0';
			when others =>
				save <= '0';
				init <= '0';
				done <= '0';
		end case;
	end process signals_gen;

	x_mux : process(x0, x_add_sub_out, init)
	begin
		if (init = '0') then
			x_mux_out <= x_add_sub_out;
		else
			x_mux_out <= x0;
		end if;
	end process x_mux;

	y_mux : process(y0, y_add_sub_out, init)
	begin
		if (init = '0') then
			y_mux_out <= y_add_sub_out;
		else
			y_mux_out <= y0;
		end if;
	end process y_mux;

	z_mux : process(angle, z_reg_out, init)
	begin
		if (init = '0') then
			z_mux_out <= z_reg_out;
		else
			z_mux_out <= angle;
		end if;
	end process z_mux;

	z_delta_mux : process(gt_hPI_s, lt_mhPI_s, init, atan_lut_out)
	begin
		if (init = '1') then
			if (gt_hPI_s = '1' or lt_mhPI_s = '1') then
				z_delta_mux_out <= HALF_PI_FX316_V;
			else
				z_delta_mux_out <= ZERO_FX316_V;
			end if;
		else
			z_delta_mux_out <= atan_lut_out;
		end if;
	end process z_delta_mux;

	z_add_sub_op_proc : process(init, z_msb, lt_mhPI_s)
	begin
		if (init = '0') then
			z_add_sub_op <= z_msb;
		else
			z_add_sub_op <= lt_mhPI_s; -- Si estoy inicializando, en funci�n de > PI/2 o < -PI/2 debo insertar como valor inicial el �ngulo original decrementado / incrementado
		end if;
	end process z_add_sub_op_proc;

	n_z_msb <= not z_msb;
end beh;
