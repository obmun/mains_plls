--------------------------------------------------------------------------------
-- *** Brief description ***
--
-- Block for managing SPI programmable ADC pre-amp (LTC 6912-1)
--
-- *** Description ***
--
-- A SPI programmable amp is found on the input stage of the ADC on the Digilent Spartan 3E board.
-- It's necessary to program this element.
--
-- This block takes care of all the digital (SPI) interfacing with the amp
--
-- ** Necessity of this block **
--
-- On initial power up (with SHDN signal open), or coming out of the hardware shutdown mode (pulling SHDN
-- to V–), both amplifiers are reset into the power-on reset state (software shutdown mode, state =
-- 8) for both channels.
--
-- En ese estado "inicial" de soft-reset, los dos amplificadores están _deshabilitados_ (entradas a
-- tercer estado)
--
-- ** The prog amp interface **
--
-- Se carga MSB first con 8 bits de datos:
-- [Q7 | Q6 | Q5 | Q4 | Q3 | Q2 | Q1 | Q0]
-- Q7 a Q4 (nibble superior) son la ganancia del canal B
-- Q3 a Q0 (nibble inferior) son la ganancia del canal A
--
-- ** Ports description **
--
-- Control and interfacing ports:
-- 1) clk: main input clock. Entity expects a hardcoded clock freq of 12.5 MHz. Block works at clk
-- rising edge
-- 2) rst: async reset
-- 3) a_gain: 4 bits for A channel gain. Used when a gain programming order (set_gain port) is executed
-- 4) b_gain: 4 bits for B channel gain. Used when a gain programming order (set_gain port) is executed
-- 5) set_gain: port similar to the "run" port of a run_done iface, which launches a gain
-- programming order. When started, done port goes down inmediately. The cycle before the operation
-- is completely finished, port goes high again.
--
-- SPI related ports
-- 1) spi_mosi: the output data generated for the amp (which should go into amp DIN pin)
-- 2) spi_sck: SPI clock output
-- 3) spi_miso: the data generated by the amp (on its DOUT pin)
-- 4) amp_ncs: the negated CS signal for the amp (pin nCS/LD on the IC)

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use WORK.COMMON.ALL;

entity prog_amp is
     port (
          clk : in std_logic;
          rst : in std_logic;
          a_gain, b_gain : in std_logic_vector(3 downto 0);
          set_gain : in std_logic;
          done: out std_logic;
          spi_owned_out : out std_logic;
          spi_mosi, spi_sck : out std_logic;
          spi_miso          : in  std_logic;
          amp_ncs           : out std_logic);
end entity prog_amp;


architecture beh of prog_amp is
     -- Global state
     type global_state_t is (
	  GLOBAL_ST_IDLE, GLOBAL_ST_GAIN_PROG);
     
     signal global_st : global_state_t;

     -- Gain programming state
     type gain_prog_state_t is (
	  GP_ST_STOPPED, GP_ST_RUNNING, GP_ST_LAST);
     
     signal gp_st : gain_prog_state_t;

     constant GP_CTR_SIZE : natural := 3;
     constant GAIN_DATA_SIZE : natural := 8;  -- Two gain registers, 4 bits each. Total: 8 bits
     
     -- Gain programming signals
     signal run_gain_prog_s, gain_prog_done_s : std_logic;
     
     signal gp_cnt : std_logic_vector(GP_CTR_SIZE - 1 downto 0); -- 3 bit counter
     signal gp_ctr_reset_s : std_logic;

     signal gain_data_reg_load_s, gp_data_MSB_s : std_logic;

     signal amp_ncs_GP_s, spi_mosi_GP_s : std_logic;
     signal enable_spi_clk_GP_s, force_high_spi_clk_GP_s : std_logic;

     signal garbage_s : std_logic_vector(GAIN_DATA_SIZE - 2 downto 0);
begin
     
     global_state_ctrl : process(clk, rst, set_gain, gain_prog_done_s)
     begin
	  if (rst = '1') then
	       global_st <= GLOBAL_ST_IDLE;
	  else
	       if (rising_edge(clk)) then
		    case global_st is
			 when GLOBAL_ST_IDLE =>
			      if (set_gain = '1') then
				   global_st <= GLOBAL_ST_GAIN_PROG;
			      else
				   global_st <= GLOBAL_ST_IDLE;
			      end if;
			 when GLOBAL_ST_GAIN_PROG =>
                              if (gain_prog_done_s = '1') then
                                   global_st <= GLOBAL_ST_IDLE;
                              else
                                   global_st <= GLOBAL_ST_GAIN_PROG;
                              end if;
			 when others =>
			      global_st <= global_st;
			      report "Unknown global state! Should not happen!" severity error;
		    end case;
	       end if;
	  end if;
     end process global_state_ctrl;

     -- Takes care of:
     -- External signals:
     -- spi_owned_out
     -- done
     -- 
     global_signal : process(global_st, gain_prog_done_s, set_gain)
     begin
	  case global_st is
	       when GLOBAL_ST_IDLE =>
                    -- External
                    spi_owned_out <= '0';
                    
                    done <= '1';

                    -- Internal
                    run_gain_prog_s <= set_gain;
	       when GLOBAL_ST_GAIN_PROG =>
                    spi_owned_out <= '1';
                    
                    done <= gain_prog_done_s;

                    -- Internal
                    run_gain_prog_s <= '0';
	       when others =>
                    spi_owned_out <= '0';

                    done <= '1';

                    -- Internal
                    run_gain_prog_s <= '0';

                    report "Unknown global state!!! Should not happen!!!"
			 severity error;
	  end case;
     end process;

     -- Gain programming state control
     gp_state_ctrl : process(clk, rst, run_gain_prog_s)
     begin
	  if (rst = '1') then
	       gp_st <= GP_ST_STOPPED;
	  else
	       if (rising_edge(clk)) then
		    case gp_st is
			 when GP_ST_STOPPED =>
			      if (run_gain_prog_s = '1') then
				   gp_st <= GP_ST_RUNNING;
			      else
				   gp_st <= GP_ST_STOPPED;
			      end if;
			 when GP_ST_RUNNING =>
                              -- This is already the _LAST_ bit, but ...
                              -- On _current_ cycle, I set the current data bit, but bit is not
                              -- stored by the amp until rising edge of beggining of next cycle.
                              -- So, I need a LAST cycle just for the final rising edge, nothing more.
                              if (to_integer(unsigned(gp_cnt)) = 7) then
                                   gp_st <= GP_ST_LAST;
                              else
                                   gp_st <= GP_ST_RUNNING;
                              end if;
                         when GP_ST_LAST =>
                              gp_st <= GP_ST_STOPPED;
			 when others =>
			      gp_st <= gp_st;
			      report "Unknown gain programming state! Should not happen!"
                                   severity error;
		    end case;
	       end if;
	  end if;
     end process;

     
     gain_programming_signals : process(gp_st, run_gain_prog_s)
     begin
          case gp_st is
	       when GP_ST_STOPPED =>
                    gain_prog_done_s <= '1';

                    -- Internal signals
                    gp_ctr_reset_s <= '1';
                    gain_data_reg_load_s <= run_gain_prog_s;

                    enable_spi_clk_GP_s <= '0';
                    force_high_spi_clk_GP_s <= '0';
                    
                    -- External signals
                    amp_ncs_GP_s <= '1';
	       when GP_ST_RUNNING =>
                    gain_prog_done_s <= '0';

                    -- Internal signals
                    gp_ctr_reset_s <= '0';
                    gain_data_reg_load_s <= '0';

                    enable_spi_clk_GP_s <= '1';
                    force_high_spi_clk_GP_s <= '0';

                    -- External signals
                    amp_ncs_GP_s <= '0';  -- Enable the device
               when GP_ST_LAST =>
                    gain_prog_done_s <= '1';

                    -- Internal signals
                    gp_ctr_reset_s <= '0';
                    gain_data_reg_load_s <= '0';

                    enable_spi_clk_GP_s <= '1';
                    force_high_spi_clk_GP_s <= '1';

                    -- External signals
                    amp_ncs_GP_s <= '0';  -- We must make sure the last rising edge (the one at the
                                          -- begging of this cycle) goes in

	       when others =>
                    report "Unknown gain programming state! Should not happen!"
			 severity error;
	  end case;
     end process;     

     -- Takes care of the gain programming counter (3 bits)
     --
     -- The gain programming counter counts from 0 to 7, counting the bits which must be send to the
     -- programmable amp.
     --
     -- Every functionality is sync.
     -- Has:
     -- * Reset (sets counter to 0)
     -- Doesn't have:
     -- * Enable. If clocked, 
     -- Outputs: dac_cnt
     gp_ctr : process(clk, gp_ctr_reset_s)
     begin
	  if (rising_edge(clk)) then
               if (gp_ctr_reset_s = '1') then
                    gp_cnt <= std_logic_vector(to_unsigned(0, GP_CTR_SIZE));
               else
                    if (to_integer(unsigned(gp_cnt)) = (2**GP_CTR_SIZE - 1)) then
                         gp_cnt <= std_logic_vector(to_unsigned(0, GP_CTR_SIZE));
                    else
                         gp_cnt <= std_logic_vector(to_unsigned(to_integer(unsigned(gp_cnt)) + 1, GP_CTR_SIZE));
                    end if;
               end if;
	  end if;
     end process;

     gain_data_reg : entity work.shift_reg(alg)
          generic map (
               width => GAIN_DATA_SIZE,
               dir => SD_LEFT,          -- According to LTC datasheet, data is MSB first
               step_s => 1)
          port map (
               clk => clk,
               load => gain_data_reg_load_s,
               we => '1',
               s_in => (others => '0'),             -- It doesn't mind the real value
               p_in(3 downto 0) => a_gain,
               p_in(GAIN_DATA_SIZE - 1 downto 4) => b_gain,
               o(GAIN_DATA_SIZE - 2 downto 0) => garbage_s,
               o(GAIN_DATA_SIZE - 1) => gp_data_MSB_s);
     spi_mosi_GP_s <= gp_data_MSB_s;

     amp_ncs <= amp_ncs_GP_s;
     spi_mosi <= spi_mosi_GP_s;
     spi_sck <= (clk and enable_spi_clk_GP_s) or force_high_spi_clk_GP_s;
end architecture beh;
