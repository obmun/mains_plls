--------------------------------------------------------------------------------
-- Company: UVigo
-- Engineer: Jacobo Cabaleiro
--
-- Create Date:    
-- Design Name:    
-- Module Name:    cordic - beh
-- Project Name:   
-- Target Device:  
-- Tool versions:  
--
-- === SPECS ===
-- Latency: VARIABLE (depends on pipeline precision)
-- Throughoutput: VARIABLE (depends on pipeline precision)
-- 
-- === Brief DESCRIPTION ===
-- Cordic based sequential engine for generating sin and cosine values from radian 
-- angles.
-- 
-- === Description ===
-- Sequential iterative cordic based sin / cos calculator. Works on clock
-- rising edge and includes a synchronous reset signal so it can be put on a known
-- state (done state).
--
-- == # of iterations ==
-- Iterations are runned till max prec on remainder angle or cos / sin value is achieved.
-- What is this limit?
-- We know on each iteration we have to possible limiting prec operations:
-- * Multiplicacion of x / y register by the correct angle (SHIFT operation),
-- for its later addition / substraction.
-- * Addition / substraction of the correspondent angle to the z register
-- (remainder angle).
-- When ANY of the previous operations reaches a precision limit, Cordic
-- algorithm must be stopped.
--
-- = Precision on shift operation =
-- On step n, precision for shift operation is n.
-- First angle (45�) starts with a tan value of 1. Consecutive angles need 1
-- more bit precsion (2^-n).
-- The problem IS ... multiplication operation!!!! COMPLETE ME!!
-- Precision on the add operation is the same: prec. on the pipeline.
-- Therefore, on the cos / sin calc, **for n prec bits, n max steps are possible**.
-- 
-- = Precision on remainder angle calc =
-- The prec on this operation is impossed by the angle values for the given
-- step / atan value, stored in the LUT. From an study of the angle values, it
-- can be clearly seen that:
-- * Every used angle is < 1 (45 � in rads is < 1) => we need a least 1 bit prec
-- even for the 1st step
-- * In the complete table, each angle requires at least 1 more prec bit than
-- previous value. THERE is one exception to this rule: rounding makes that 7th
-- and 8th angles msb is the same. Ignoring this anomality, we can MAKE THE FOLLOWING RULE: for each
-- step, angle needs 1 more bit of prec.
--
-- Therefore, **if we have n bits prec, at most n different angles can be added / subs
-- from z**.
--
-- Both restrictions are EQUIVALENT [but remember, we have the exception to the
-- precision on remainder angle] => *for n prec bits, max n steps can be run*.
-- 
-- == Ports ==
-- * Inputs *
-- -> CLK
-- -> RST: synchronous reset
-- -> RUN: run/done iface run signal. See below for description
-- -> ANGLE: input angle, in radians
-- * Outputs *
-- -> SIN: sin value for given input angle
-- -> COS: cos value for given input angle
-- -> DONE: run/done iface done signal. See below for description
--
-- Dependencies:
-- 
-- === Changelog ===
-- Revision 0.04 - Made parametrizable.
-- MARK -> revision 0.03 has been tested. Works OK. Small problems with
-- precision appear near 0 radians
-- Revision 0.03 - Counter reset is now synchronous (UNTESTED)
-- Revision 0.02 - New state machine (TESTED)
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use WORK.COMMON.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.all;

entity cordic is
        -- rev 0.04
	generic (
		width : natural := PIPELINE_WIDTH;
                prec : natural := PIPELINE_PREC);
	port (
		clk, rst, run : in std_logic;
		angle : in std_logic_vector(width - 1 downto 0); -- In RADIANS!
		sin, cos : out std_logic_vector(width - 1 downto 0);
		done : out std_logic);
end cordic;

architecture beh of cordic is
	type state_t is (
		ST_DONE, ST_INIT, ST_RUNNING, ST_LAST
	);

	signal st : state_t; -- Se podr�a hacer con una variable compartida, aunque debido al posible comportamiento no determinista se prefiere simular (como en la realidad) mediante una se�al
        
	signal step : natural;

	-- Control signas (generated by FSM)
	signal init, save : std_logic;

	-- Cordic interconnect signals
	signal x0, y0 : std_logic_vector(width - 1 downto 0);
	signal gt_hPI_s, lt_mhPI_s : std_logic;
	signal z_add_sub_op : std_logic;
	signal x_mux_out, y_mux_out, z_mux_out : std_logic_vector(width - 1 downto 0);
	signal z_delta_mux_out, atan_lut_out : std_logic_vector(width - 1 downto 0);
	signal x_reg_out, y_reg_out, z_reg_out : std_logic_vector(width - 1 downto 0);
	signal x_add_sub_out, y_add_sub_out, z_add_sub_out : std_logic_vector(width - 1 downto 0);
	signal x_shift_out, y_shift_out : std_logic_vector(width - 1 downto 0);

	alias z_msb : std_logic is z_reg_out(width - 1);
	signal n_z_msb : std_logic;

	-- Components
	component add_sub is
		generic (
			width : natural := PIPELINE_WIDTH
		);
		port (
			a, b: in std_logic_vector(width - 1 downto 0);
			add_nsub : in std_logic;
			o: out std_logic_vector(width - 1 downto 0);
			f_ov, f_z: out std_logic
		);
	end component;

	component reg is
		generic (
			width : natural := PIPELINE_WIDTH
		);
		port (
			clk, we, rst : in std_logic;
			i : in std_logic_vector (width - 1 downto 0);
			o : out std_logic_vector (width - 1 downto 0)
		);
	end component;

	component k_lt_comp is
		generic (
			width : natural := PIPELINE_WIDTH;
			k : pipeline_integer := 0
		);
		port (
			a : in std_logic_vector(width - 1 downto 0);
			a_lt_k : out std_logic
		);
	end component;

	component k_gt_comp is
		generic (
			width : natural := PIPELINE_WIDTH;
			k : pipeline_integer := 0
		);
		port (
			a : in std_logic_vector(width - 1 downto 0);
			a_gt_k : out std_logic
		);
	end component;

begin
        -- Is input angle < - PI / 2.0?
	lt_comp : k_lt_comp
		generic map (
                        width => width,
			k => to_integer(MINUS_HALF_PI, width, prec))
		port map (
			a => angle,
			a_lt_k => lt_mhPI_s);

        -- Is input angle > PI / 2.0?
	gt_comp : k_gt_comp
		generic map (
                        width => width, 
			k => to_integer(HALF_PI, width, prec))
		port map (
			a => angle,
			a_gt_k => gt_hPI_s);

	x_add_sub : add_sub
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => x_reg_out,
			b => y_shift_out,
			add_nsub => z_msb,
			-- SALIDAS
			o => x_add_sub_out,
                        -- Unconnected
                        f_ov => open,
                        f_z => open);

	y_add_sub : add_sub
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => y_reg_out,
			b => x_shift_out,
			add_nsub => n_z_msb,
			-- SALIDAS
			o => y_add_sub_out,
                        -- Unconnected
                        f_ov => open,
                        f_z => open);

	z_add_sub : add_sub
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => z_mux_out,
			b => z_delta_mux_out,
			add_nsub => z_add_sub_op,
			-- SALIDS
			o => z_add_sub_out);

	x_reg : reg
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => x_mux_out,
			-- SALIDAS
			o => x_reg_out);

	y_reg : reg
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => y_mux_out,
			-- SALIDAS
			o => y_reg_out);

	z_reg : reg
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => z_add_sub_out,
			-- SALIDAS
			o => z_reg_out);

        -- Final cos value storage. Does not take an active part in algorithm
	cos_reg : reg
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => save, rst => rst,
			i => x_add_sub_out,
			-- SALIDAS
			o => cos);

        -- Final sin value storage. Does not take an active part in algorithm
	sin_reg : reg
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => save, rst => rst,
			i => y_add_sub_out,
			-- SALIDAS
			o => sin);

	x_shifter : entity work.signed_r_shifter(beh)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			i => x_reg_out,
			n => step,
			-- SALIDAS
			o => x_shift_out);

	y_shifter : entity work.signed_r_shifter(beh)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			i => y_reg_out,
			n => step,
			-- SALIDAS
			o => y_shift_out);

	atan_lut : entity work.cordic_atan_lut(beh)
                generic map (
                        width      => width,
                        prec       => prec,
                        last_angle => prec - 1)
		port map (
			addr  => step,
			angle => atan_lut_out);

	n_z_msb <= not z_msb;

        -- ********************************************
        -- * Componentes for ALGORITHM initialization *
        -- ********************************************
        -- Mux for x reg input. Allows correct initialization of x during init.
	x_mux : process(x0, x_add_sub_out, init)
	begin
		if (init = '0') then
			x_mux_out <= x_add_sub_out;
		else
			x_mux_out <= x0;
		end if;
	end process x_mux;

                -- Mux for y reg input. Same function as x reg but for y reg.
	y_mux : process(y0, y_add_sub_out, init)
	begin
		if (init = '0') then
			y_mux_out <= y_add_sub_out;
		else
			y_mux_out <= y0;
		end if;
	end process y_mux;

        -- Initialization of the z (angle) register
	z_mux : process(angle, z_reg_out, init)
	begin
		if (init = '0') then
			z_mux_out <= z_reg_out;
		else
			z_mux_out <= angle;
		end if;
	end process z_mux;

        -- Sets a special initial value for the 2nd operand of the z reg adder
	z_delta_mux : process(gt_hPI_s, lt_mhPI_s, init, atan_lut_out)
	begin
		if (init = '1') then
			if (gt_hPI_s = '1' or lt_mhPI_s = '1') then
				z_delta_mux_out <= to_vector(HALF_PI, width, prec);
			else
				z_delta_mux_out <= (others => '0');
			end if;
		else
			z_delta_mux_out <= atan_lut_out;
		end if;
	end process z_delta_mux;
        
        -- Process which takes care of selecting the correct init values for x and
        -- y registers depending on the quadrant of the input angle
	cordic_elem_init : process(gt_hPI_s, lt_mhPI_s)
	begin
		if (gt_hPI_s = '1') then
			x0 <= (others => '0');
			y0 <= to_vector(INV_CORDIC_GAIN, width, prec);
		elsif (lt_mhPI_s = '1') then
			x0 <= (others => '0');
			y0 <= to_vector(MINUS_INV_CORDIC_GAIN, width, prec);
		else
			x0 <= to_vector(INV_CORDIC_GAIN, width, prec);
			y0 <= (others => '0');
		end if;
	end process;

        z_add_sub_op_proc : process(init, z_msb, lt_mhPI_s)
	begin
		if (init = '0') then
			z_add_sub_op <= z_msb;
		else
			z_add_sub_op <= lt_mhPI_s; -- Si estoy inicializando, en funci�n de > PI/2 o < -PI/2 debo insertar como valor inicial el �ngulo original decrementado / incrementado
		end if;
	end process z_add_sub_op_proc;

        
        -- *******************
        -- * State processes *
        -- *******************
        
        -- Counter process. For the internal process counter.
        -- # of steps = PREC BITS! See description for more info
	step_counter : process(clk)
		variable step_counter : std_logic_vector((integer(round(ceil(log2(real(prec - 1))))) - 1) downto 0);
	begin
                assert false report "Cordic step counter width: " & integer'image(integer(round(ceil(log2(real(prec)))))) severity note;
                
		if (rising_edge(clk)) then
			if (init = '1') then
				step_counter := (others => '0');
			else
                                -- To achieve an OPTIMAL counter size, make it
                                -- fold the CORRECT WAY (on saturation of
                                -- optimun width)
                                if (unsigned(step_counter) = (integer(round(2.0 ** ceil(log2(real(prec - 1))))) - 1)) then
                                        step_counter := (others => '0');
                                else
                                        step_counter := std_logic_vector(unsigned(step_counter) + 1);
                                end if;
			end if;
		end if;
		step <= to_integer(unsigned(step_counter));
	end process;


        state_ctrl : process(clk, run, rst)
	begin
		if (rising_edge(clk)) then
			if (rst = '1') then
				st <= ST_DONE;
			else
				case st is
					when ST_DONE =>
						if (run = '1') then
							st <= ST_INIT;
						else
							st <= ST_DONE;
						end if;
					when ST_INIT =>
						st <= ST_RUNNING;
					when ST_RUNNING =>
						if (step = prec - 1) then
							st <= ST_LAST;
						else
							st <= ST_RUNNING;
						end if;
					when ST_LAST =>
                                                st <= ST_DONE;
					when others =>
						assert false
							report "Unkown Cordic state! Should not happen!"
							severity error;
						st <= st;
				end case;
			end if;
		end if;
	end process state_ctrl;

	signals_gen : process(st)
	begin
		case st is
			when ST_DONE =>
				init <= '0';
				save <= '0';
				done <= '1';
			when ST_INIT =>
				init <= '1';
				save <= '0';
				done <= '0';
			when ST_RUNNING =>
				init <= '0';
				save <= '0';
				done <= '0';
			when ST_LAST =>
				save <= '1';
				init <= '0';
				done <= '0';
			when others =>
				save <= '0';
				init <= '0';
				done <= '0';
		end case;
	end process signals_gen;
end beh;
