--------------------------------------------------------------------------------
-- Company: UVigo
-- Engineer: Jacobo Cabaleiro
--
-- Create Date:    
-- Design Name:    
-- Module Name:    fa - beh
-- Project Name:  
-- Target Device:  
-- Tool versions: 
--
-- *** SPECS ***
-- Latency: 1 clk [when waken up] / 0 clks
-- Troughoutput: 1 sample / cycle
-- 
-- *** BRIEF DESCRIPTION ***
-- Class: sequential
-- Moving Averega Filter, recursive implementation, with configurable delay (rejected harmonic frequencies thru generic ports.
-- Works on clock's rising edge and has synchronous reset.
-- 
-- *** DESCRIPTION ***
-- Includes a synchronous reset.
-- It's an IIR, so you should be using a LOT OF PRECISION!!! when implementing
-- this thing. You have been warned.
-- 
-- == PORT DESCRIPTION ==
-- = Generics =
-- * width: ports and internal pipeline width
-- * prec: ports and internal pipeline precision
-- * delay: # of clocks of delay (at least 1)
-- 
-- *** Changelog ***
-- Revision 0.05 - Stop fucking, please. CHANGED the implementation. This is
-- the REAL ONE. Check PFC notes.
-- Revision 0.04 - With change of kcm, no input multiplying constant is real
-- and user must not scale it by SAMPLING_PERIOD as its done inside the kcm_integrator.
-- Revision 0.03 - Implement new seq. control iface. REALLY create the generic
-- for freq. and k control, instead of just advertising it in the brief description
-- Revision 0.02 - Added run / done style PORTS for syncronization with other sequential algorithms.
-- Revision 0.01 - File Created
--
-- *** Todo ***
-- | 1.- REVIEW SINTHESIS!!!
-- | 2.- Correctly implement RST behaviour!!!
--------------------------------------------------------------------------------

library IEEE;
library WORK;
use WORK.COMMON.all;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity fa is
        -- rev 0.04
        generic (
                width : natural := PIPELINE_WIDTH;
                prec : natural := PIPELINE_PREC;
                delay : natural; 
                -- Seq. block iface
                delayer_width : natural := 1);
	port (
		clk, rst : in std_logic;
		i : in std_logic_vector(width - 1 downto 0);
		o : out std_logic_vector(width - 1 downto 0);
                run_en : in std_logic;
                run_passthru : out std_logic;
                delayer_in : in std_logic_vector(delayer_width - 1 downto 0);
                delayer_out : out std_logic_vector(delayer_width - 1 downto 0));
end fa;

architecture beh of fa is
        constant d_inv : real := 1.0 / real(delay);
	signal kcm_out_s, fifo_out_s, reg_out_s, sub_out_s, o_s : std_logic_vector(width - 1 downto 0);
        signal delayer_in_s, delayer_out_s : std_logic_vector(delayer_width - 1 downto 0);        
begin
        kcm_i : entity work.kcm(beh)
                generic map (
                        width => width,
                        prec  => prec,
                        k     => d_inv)
                port map (
                        i => i,
                        o => kcm_out_s);

	fifo_i : entity work.fifo(alg)
		generic map (
                        width => width,
                        size => delay)
		port map (
			i => kcm_out_s,
			o => fifo_out_s,
			clk => clk, we => run_en);

	sub_i : entity work.subsor(alg)
		generic map (
                        width => width)
		port map (
			a => kcm_out_s,
			b => fifo_out_s,
			o => sub_out_s,
                        -- Unconnected
                        f_ov => open,
                        f_z => open);

        reg_i : entity work.reg(alg)
                generic map (
                        width => width)
                port map (
                        clk => clk,
                        we  => run_en,
                        rst => rst,
                        i   => o_s,
                        o   => reg_out_s);

        add_i : entity work.adder(alg)
                generic map (
                        width => width)
                port map (
                        a    => sub_out_s,
                        b    => reg_out_s,
                        o    => o_s,
                        f_ov => open,
                        f_z  => open);

        o <= o_s;

        delayer : entity work.reg(alg)
                generic map (
                        width => delayer_width)
		port map (
			clk => clk, we => '1', rst => rst,
			i => delayer_in_s,
			o => delayer_out_s);

        single_delayer_gen: if (delayer_width = 1) generate
                delayer_in_s(0) <= run_en;
                run_passthru <= std_logic(delayer_out_s(0));
                delayer_out(0) <= delayer_out_s(0);
        end generate single_delayer_gen;
        
        broad_delayer_gen: if (delayer_width > 1) generate
                delayer_in_s(0) <= run_en;
                delayer_in_s(delayer_width - 1 downto 1) <= delayer_in(delayer_width - 1 downto 1);
                run_passthru <= std_logic(delayer_out_s(0));
                delayer_out <= delayer_out_s;
        end generate broad_delayer_gen;
end beh;
