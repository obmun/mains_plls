--------------------------------------------------------------------------------
-- Company: UVigo
-- Engineer: Jacobo Cabaleiro
--
-- Create Date:    
-- Design Name:    
-- Module Name:    cordic - beh
-- Project Name:   
-- Target Device:  
-- Tool versions:  
--
-- === SPECS ===
-- Latency: VARIABLE (depends on pipeline precision)
-- Throughoutput: VARIABLE (depends on pipeline precision)
-- 
-- === Brief DESCRIPTION ===
-- Cordic based sequential engine for calculating atan2 and hypot (vector modulus).
-- Based on a CORDIC engine working in vectoring mode
-- 
-- === Description ===
--
-- == # of iterations ==
-- See cordic.vhd
--
-- == Ports ==
-- * Inputs *
-- -> CLK
-- -> RST: synchronous reset
-- -> RUN: run/done iface run signal. See block_interfaces.txt for description
-- -> X:
-- -> Y:
-- * Outputs *
-- -> ANGLE:
-- -> MOD:
-- -> DONE: run/done iface done signal. See below for description
--
-- Dependencies:
-- 
-- === Changelog ===
-- Revision 0.01 - File created, based on cordic.vhd
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use WORK.COMMON.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.all;

entity cordic_atan is
        -- rev 0.01
	generic (
		width : natural := PIPELINE_WIDTH;
                prec : natural := PIPELINE_PREC);
	port (
		clk, rst, run : in std_logic;
		x, y : in std_logic_vector(width - 1 downto 0);
		angle, modu : out std_logic_vector(width - 1 downto 0);
		done : out std_logic);
end cordic_atan;

architecture structural of cordic_atan is
	type state_t is (
		ST_DONE, ST_INIT, ST_RUNNING, ST_LAST
	);

	signal st : state_t; -- Se podr�a hacer con una variable compartida, aunque debido al posible comportamiento no determinista se prefiere simular (como en la realidad) mediante una se�al
        
	signal step_s : natural;

	-- Control signals (generated by FSM)
	signal init_s, save_s : std_logic;

	-- Cordic interconnect signals
	signal x0_s, y0_s, z0_s : std_logic_vector(width - 1 downto 0);
	signal x_lt_0_s, y_lt_0_s : std_logic;
	signal z_add_sub_op_s : std_logic;
	signal x_mux_out_s, y_mux_out_s, z_mux_out_s : std_logic_vector(width - 1 downto 0);
	signal atan_lut_out_s : std_logic_vector(width - 1 downto 0);
	signal x_reg_out_s, y_reg_out_s, z_reg_out_s : std_logic_vector(width - 1 downto 0);
	signal x_add_sub_out_s, y_add_sub_out_s, z_add_sub_out_s : std_logic_vector(width - 1 downto 0);
        signal modu_reg_out_s : std_logic_vector(width - 1 downto 0);
	signal x_shift_out_s, y_shift_out_s : std_logic_vector(width - 1 downto 0);

	alias y_msb_s : std_logic is y_reg_out_s(width - 1);
	signal n_y_msb_s : std_logic;

        pure function cordic_gain ( n_iters : natural ) return real is
                variable tmp_gain : real := 1.0;
        begin
                for i in 0 to n_iters - 1 loop
                        tmp_gain := tmp_gain * sqrt(1.0 + 2.0 ** (-2.0 * real(i)));
                end loop;
                return tmp_gain;
        end;
begin
        -- Is x input < 0?
        x_lt_0_s <= x(width - 1);
        -- Is y input < 0?
        y_lt_0_s <= y(width - 1);
        
	x_add_sub : entity work.add_sub(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => x_reg_out_s,
			b => y_shift_out_s,
			add_nsub => n_y_msb_s,
			-- SALIDAS
			o => x_add_sub_out_s,
                        -- Unconnected
                        f_ov => open,
                        f_z => open);

	y_add_sub : entity work.add_sub(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => y_reg_out_s,
			b => x_shift_out_s,
			add_nsub => y_msb_s,
			-- SALIDAS
			o => y_add_sub_out_s,
                        -- Unconnected
                        f_ov => open,
                        f_z => open);

	z_add_sub : entity work.add_sub(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			a => z_reg_out_s,
			b => atan_lut_out_s,
			add_nsub => z_add_sub_op_s,
			-- SALIDS
			o => z_add_sub_out_s);

	x_reg : entity work.reg(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => x_mux_out_s,
			-- SALIDAS
			o => x_reg_out_s);

	y_reg : entity work.reg(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => y_mux_out_s,
			-- SALIDAS
			o => y_reg_out_s);

        n_y_msb_s <= not y_msb_s;

	z_reg : entity work.reg(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => '1', rst => '0',
			i => z_mux_out_s,
			-- SALIDAS
			o => z_reg_out_s);

        -- Final vector modulus value storage. It's not an active part of the algorithm

        
	modu_reg : entity work.reg(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => save_s, rst => rst,
			i => x_add_sub_out_s,
			-- SALIDAS
			o => modu_reg_out_s);

        modu_kcm : entity work.kcm(structural_mm)
                generic map (
                        width => width,
                        prec  => prec,
                        k     => 1.0/cordic_gain(prec))
                port map (
                        i => modu_reg_out_s,
                        o => modu);

        -- Final vector phase (atan2) value storage. It's not an active part
        -- of the algorithm
	angle_reg : entity work.reg(alg)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			clk => clk, we => save_s, rst => rst,
			i => z_add_sub_out_s,
			-- SALIDAS
			o => angle);

	x_shifter : entity work.signed_r_shifter(beh)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			i => x_reg_out_s,
			n => step_s,
			-- SALIDAS
			o => x_shift_out_s);

	y_shifter : entity work.signed_r_shifter(beh)
                generic map (
                        width => width)
		port map (
			-- ENTRADAS
			i => y_reg_out_s,
			n => step_s,
			-- SALIDAS
			o => y_shift_out_s);

	atan_lut : entity work.cordic_atan_lut(beh)
                generic map (
                        width      => width,
                        prec       => prec,
                        last_angle => prec - 1)
		port map (
			addr  => step_s,
			angle => atan_lut_out_s);

        -- ********************************************
        -- * Componentes for ALGORITHM initialization *
        -- ********************************************
        -- Mux for x reg input. Allows correct initialization of x during init.
	x_mux : process(x0_s, x_add_sub_out_s, init_s)
	begin
		if (init_s = '0') then
			x_mux_out_s <= x_add_sub_out_s;
		else
			x_mux_out_s <= x0_s;
		end if;
	end process x_mux;

                -- Mux for y reg input. Same function as x reg but for y reg.
	y_mux : process(y0_s, y_add_sub_out_s, init_s)
	begin
		if (init_s = '0') then
			y_mux_out_s <= y_add_sub_out_s;
		else
			y_mux_out_s <= y0_s;
		end if;
	end process y_mux;

        -- Initialization of the z (angle) register
	z_mux : process(init_s, z_add_sub_out_s, z0_s)
	begin
		if (init_s = '0') then
			z_mux_out_s <= z_add_sub_out_s;
		else
                        z_mux_out_s <= z0_s;
		end if;
	end process z_mux;

        -- Process which takes care of selecting the correct init values for x
        -- , y, and z registers depending on the quadrant of the input vector
	cordic_elem_init : process(x_lt_0_s, y_lt_0_s, x, y)
	begin
                if (x_lt_0_s = '1') then
                        x0_s <= std_logic_vector(-signed(x));
                        y0_s <= std_logic_vector(-signed(y));
                        if (y_lt_0_s = '1') then
                                z0_s <= to_vector(MINUS_PI, width, prec);
                        else
                                z0_s <= to_vector(PI, width, prec);
                        end if;
                else
                        x0_s <= x;
                        y0_s <= y;
                        z0_s <= (others => '0');
                end if;
	end process;

        z_add_sub_op_s <= n_y_msb_s;

        
        -- *******************
        -- * State processes *
        -- *******************
        
        -- Counter process. For the internal process counter.
        -- # of steps = PREC BITS! See description for more info
	step_counter : process(clk)
		variable step_counter : std_logic_vector((integer(round(ceil(log2(real(prec - 1))))) - 1) downto 0);
	begin
                assert false report "Cordic step counter width: " & integer'image(integer(round(ceil(log2(real(prec)))))) severity note;
                
		if (rising_edge(clk)) then
			if (init_s = '1') then
				step_counter := (others => '0');
			else
                                -- To achieve an OPTIMAL counter size, make it
                                -- fold the CORRECT WAY (on saturation of
                                -- optimun width)
                                if (unsigned(step_counter) = (integer(round(2.0 ** ceil(log2(real(prec - 1))))) - 1)) then
                                        step_counter := (others => '0');
                                else
                                        step_counter := std_logic_vector(unsigned(step_counter) + 1);
                                end if;
			end if;
		end if;
		step_s <= to_integer(unsigned(step_counter));
	end process;


        state_ctrl : process(clk)
	begin
		if (rising_edge(clk)) then
			if (rst = '1') then
				st <= ST_DONE;
			else
				case st is
					when ST_DONE =>
						if (run = '1') then
							st <= ST_INIT;
						else
							st <= ST_DONE;
						end if;
					when ST_INIT =>
						st <= ST_RUNNING;
					when ST_RUNNING =>
						if (step_s = prec - 1) then
							st <= ST_LAST;
						else
							st <= ST_RUNNING;
						end if;
					when ST_LAST =>
                                                st <= ST_DONE;
					when others =>
						assert false
							report "Unkown Cordic state! Should not happen!"
							severity error;
						st <= st;
				end case;
			end if;
		end if;
	end process state_ctrl;

	signals_gen : process(st)
	begin
		case st is
			when ST_DONE =>
				init_s <= '0';
				save_s <= '0';
				done <= '1';
			when ST_INIT =>
				init_s <= '1';
				save_s <= '0';
				done <= '0';
			when ST_RUNNING =>
				init_s <= '0';
				save_s <= '0';
				done <= '0';
			when ST_LAST =>
				save_s <= '1';
				init_s <= '0';
				done <= '0';
			when others =>
				save_s <= '0';
				init_s <= '0';
				done <= '0';
		end case;
	end process signals_gen;
end structural;
