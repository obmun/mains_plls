--------------------------------------------------------------------------------
-- *** Brief description ***
-- 
-- SyncMVA synchronization scheme entity.
--
-- *** Revisions ***
--
-- - For new revision information, check Mercurial project repo
--
-- - Revision 0.01 - File Created
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.common.all;

entity p2_sync is
     port (
          clk, sample, rst : in std_logic;
          in_signal : in std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
          phase, out_signal, ampl : out std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
          done : out std_logic);
end p2_sync;

architecture structural of p2_sync is
     constant FA_PREC : natural := EXT_IIR_FILTERS_PREC;
     
     signal first_run_s, first_run_pulsed_s, freq2phase_delayed_run_s : std_logic;
     signal sincos_cordic_done_s, sincos_cordic_done_pulsed_s, sin_fa_delayed_run_s, cos_fa_delayed_run_s, fa_delayed_run_s : std_logic;
     signal atan_cordic_done_s, atan_has_run_since_sample_s : std_logic;

     signal in_signal_reg_out_s, freq2phase_out_s, freq2phase_out_REG_s, sin_s, cos_s : std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
     signal in_sin_mul_out_s, in_sin_doubler_out_s, in_cos_mul_out_s, in_cos_doubler_out_s : std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
     signal sin_speedup_reg_out_s : std_logic_vector(PIPELINE_WIDTH downto 0);
     signal cos_speedup_reg_out_s : std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
     signal in_sin_doubler_out_E_s, in_cos_doubler_out_E_s, sin_fa_out_E_s, cos_fa_out_E_s : std_logic_vector(EXT_PIPELINE_WIDTH - 1 downto 0);
     signal sin_fa_out_s, sin_fa_out_REG_s, cos_fa_out_s, cos_fa_out_REG_s, sin_sin_mul_out_s, cos_cos_mul_out_s : std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
     signal phase_error_s, big_phase_s, main_phase_det_k_s : std_logic_vector(PIPELINE_WIDTH - 1 downto 0);
begin  -- structural

     first_run_s <= atan_cordic_done_s and sample;
     first_run_pulser : entity work.done_pulser(beh)
          port map (
               clk => clk,
               en  => '1',
               rst => rst,
               i   => first_run_s,
               o   => first_run_pulsed_s);

     in_signal_reg : entity work.reg(alg)
          port map (
               clk => clk,
               we => first_run_pulsed_s,
               rst => rst,
               i => in_signal,
               o => in_signal_reg_out_s);

     -- We can't integrate a gain here, but I don't need extended precision because there is no
     -- input.
     --
     -- As every 0 latency run_passthru blocks, each time I update I generate the internal state
     -- required for the _next_ sample time. Given we have no input, the value being generated by
     -- the block before the clk pulse is already the one I need for this cycle in the rest of the
     -- elements.
     --
     -- That means run_passthru signal from this block is not needed in the rest of the
     -- elements in the case of a 0 latency block. As the signal is not delayed at all (according to
     -- the run_passthru interface specs), we can leave the CORDIC run dependant on this
     -- run_passthru output just in case in the future the impementatino of freq2phase is changed.
     --
     -- However, we need the instantaneous phase value at the final stages, so we need to register
     -- the output.
     freq2phase_i : entity work.freq2phase(beh)
          generic map (
               width         => PIPELINE_WIDTH,
               prec          => PIPELINE_PREC,
               gain          => 0.0, -- We have a 0 input. With a 0 gain we reassure that the
                                     -- input KCM on the freq2phase does not gen synthethized.
               delayer_width => 1)
          port map (
               clk => clk,
               rst => rst,
               f => to_pipeline_vector(0.0),
               p => freq2phase_out_s,
               run_en => first_run_pulsed_s,
               run_passthru => freq2phase_delayed_run_s,
               delayer_in => "-",
               delayer_out => open);

     natural_inst_phase_reg_i : entity work.reg(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               clk   => clk,
               we    => first_run_pulsed_s,
               rst   => rst,
               i     => freq2phase_out_s,
               o     => freq2phase_out_REG_s);

     sincos_cordic : entity work.cordic(structural)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               clk   => clk,
               rst   => rst,
               run   => freq2phase_delayed_run_s,
               angle => freq2phase_out_s,
               sin   => sin_s,
               cos   => cos_s,
               done  => sincos_cordic_done_s);

     sincos_cordic_done_pulser : entity work.done_pulser(beh)
          port map (
               clk => clk,
               en  => '1',
               rst => rst,
               i   => sincos_cordic_done_s,
               o   => sincos_cordic_done_pulsed_s);

     in_sin_mul : entity work.mul(beh)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               a => in_signal_reg_out_s,
               b => sin_s,
               o => in_sin_mul_out_s);

     in_sin_doubler : entity work.k_2_mul(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               i => in_sin_mul_out_s,
               o => in_sin_doubler_out_s);

     sin_speedup_reg :  entity work.reg(alg)
          generic map (
               width => PIPELINE_WIDTH + 1)
          port map (
               clk => clk,
               we => '1',
               rst => rst,
               i(PIPELINE_WIDTH - 1 downto 0) => in_sin_doubler_out_s,
               i(PIPELINE_WIDTH) => sincos_cordic_done_pulsed_s,
               o => sin_speedup_reg_out_s);

     in_cos_mul : entity work.mul(beh)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               a => in_signal_reg_out_s,
               b => cos_s,
               o => in_cos_mul_out_s);

     in_cos_doubler : entity work.k_2_mul(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               i => in_cos_mul_out_s,
               o => in_cos_doubler_out_s);

     cos_speedup_reg :  entity work.reg(alg)
          generic map (
               width => PIPELINE_WIDTH)
          -- sincos_cordic_done_pulsed_s is already delayed by sin_speedup_reg
          port map (
               clk => clk,
               we => '1',
               rst => rst,
               i => in_cos_doubler_out_s,
               o => cos_speedup_reg_out_s);

     sin_fa_input_conv : entity work.pipeline_conv(alg)
          generic map (
               in_width  => PIPELINE_WIDTH,
               in_prec   => PIPELINE_PREC,
               out_width => EXT_PIPELINE_WIDTH,
               out_prec  => FA_PREC)
          port map (
               i => sin_speedup_reg_out_s(PIPELINE_WIDTH - 1 downto 0),
               o => in_sin_doubler_out_E_s);

     -- 100 Hz tuned MVA (MAF)
     sin_fa : entity work.fa(beh)
          generic map (
               width         => EXT_PIPELINE_WIDTH,
               prec          => FA_PREC,
               delay         => 100,
               delayer_width => 1)
          port map (
               clk            => clk,
               rst            => rst,
               i              => in_sin_doubler_out_E_s,
               o              => sin_fa_out_E_s,
               run_en         => sin_speedup_reg_out_s(PIPELINE_WIDTH),
               run_passthru   => sin_fa_delayed_run_s,
               delayer_in => (others => '-'),
               delayer_out => open);
     
     sin_fa_output_conv : entity work.pipeline_conv(alg)
          generic map (
               out_width => PIPELINE_WIDTH,
               out_prec  => PIPELINE_PREC,
               in_width  => EXT_PIPELINE_WIDTH,
               in_prec   => FA_PREC)
          port map (
               i => sin_fa_out_E_s,
               o => sin_fa_out_s);

     -- FA output is direcly required (combinational) on the recovered signal output.
     -- We know that the output of this element, after the cycle it finishes calculation, is no
     -- longer valid, so it must be registered. The same happens with the cos fa output.
     sin_fa_out_reg : entity work.reg(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               clk => clk,
               we => sin_fa_delayed_run_s,
               rst => rst,
               i => sin_fa_out_s,
               o => sin_fa_out_REG_s);
     
     cos_fa_input_conv : entity work.pipeline_conv(alg)
          generic map (
               in_width  => PIPELINE_WIDTH,
               in_prec   => PIPELINE_PREC,
               out_width => EXT_PIPELINE_WIDTH,
               out_prec  => FA_PREC)
          port map (
               i => cos_speedup_reg_out_s,
               o => in_cos_doubler_out_E_s);

     cos_fa : entity work.fa(beh)
          generic map (
               width         => EXT_PIPELINE_WIDTH,
               prec          => FA_PREC,
               delay         => 100,
               delayer_width => 1)
          port map (
               clk            => clk,
               rst            => rst,
               i              => in_cos_doubler_out_E_s,
               o              => cos_fa_out_E_s,
               run_en         => sin_speedup_reg_out_s(PIPELINE_WIDTH),
               run_passthru   => cos_fa_delayed_run_s,
               delayer_in => (others => '-'),
               delayer_out => open);
     
     cos_fa_output_conv : entity work.pipeline_conv(alg)
          generic map (
               out_width => PIPELINE_WIDTH,
               out_prec  => PIPELINE_PREC,
               in_width  => EXT_PIPELINE_WIDTH,
               in_prec   => FA_PREC)
          port map (
               i => cos_fa_out_E_s,
               o => cos_fa_out_s);

     cos_fa_out_reg : entity work.reg(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               clk => clk,
               we => cos_fa_delayed_run_s,
               rst => rst,
               i => cos_fa_out_s,
               o => cos_fa_out_REG_s);

     fas_done_pulsed_and_i : entity work.pulsed_done_and(beh)
          generic map (
               width => 2)
          port map (
               clk => clk,
               rst => rst,
               i(0) => sin_fa_delayed_run_s,
               i(1) => cos_fa_delayed_run_s,
               o => fa_delayed_run_s);

     atan_cordic : entity work.cordic_atan(structural)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               clk => clk,
               rst => rst,
               run => fa_delayed_run_s,
               x => sin_fa_out_s,
               y => cos_fa_out_s,
               angle => phase_error_s,
               modu => ampl,
               done  => atan_cordic_done_s);

     -- We're using a 3 bits magn pipeline, that is we have the range (-8, 7.999), enough even for a
     -- full pi phase correction (output of the atan element is on the (-pi, pi) range).
     phase_adder : entity work.adder(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               a => phase_error_s,
               b => freq2phase_out_REG_s,
               o => big_phase_s);

     -- Phase correction
     phase_correctin: block is
     begin
          main_phase_det_k_gen : process(big_phase_s)
          begin
               if (signed(big_phase_s) > signed(to_pipeline_vector(PI))) then
                    main_phase_det_k_s <= to_pipeline_vector(MINUS_TWO_PI);
               elsif (signed(big_phase_s) < signed(to_pipeline_vector(MINUS_PI))) then
                    main_phase_det_k_s <= to_pipeline_vector(TWO_PI);
               else
                    main_phase_det_k_s <= (others => '0');
               end if;
          end process main_phase_det_k_gen;
          main_phase_det_adder : entity work.adder(alg)
               generic map (
                    width => PIPELINE_WIDTH)
               port map (
                    a => big_phase_s,
                    b => main_phase_det_k_s,
                    o => phase);          
     end block;

     -- done signal generation
     done_signal_gen: block is
     begin
          -- Some extra processes needed to make done behave according to
          -- block_interface.txt specifications
          atan_has_run_since_sample_gen : process(clk, sample, rst, fa_delayed_run_s)
          begin
               if rising_edge(clk) then
                    if (rst = '1') then
                         atan_has_run_since_sample_s <= '1';
                    else
                         if (sample = '1') then
                              atan_has_run_since_sample_s <= '0';
                         else
                              if (fa_delayed_run_s = '1') then
                                   atan_has_run_since_sample_s <= '1';
                              end if;
                         end if;
                    end if;
               end if;
          end process atan_has_run_since_sample_gen;
          -- On the switch below we generate a little glitch to one of 1 or 2 ticks on the done signal, but it's
          -- after the rising edge of clk, so it's benign.
          done <= atan_cordic_done_s when atan_has_run_since_sample_s = '1' else '0';          
     end block done_signal_gen;

     sin_sin_mul : entity work.mul(beh)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               a => sin_s,
               b => sin_fa_out_REG_s,
               o => sin_sin_mul_out_s);

     cos_cos_mul : entity work.mul(beh)
          generic map (
               width => PIPELINE_WIDTH,
               prec  => PIPELINE_PREC)
          port map (
               a => cos_s,
               b => cos_fa_out_REG_s,
               o => cos_cos_mul_out_s);

     out_signal_adder_i : entity work.adder(alg)
          generic map (
               width => PIPELINE_WIDTH)
          port map (
               a => sin_sin_mul_out_s,
               b => cos_cos_mul_out_s,
               o => out_signal);
end structural;
