--------------------------------------------------------------------------------
-- Company: Universidad de Vigo
-- Engineer: Jacobo Cabaleiro
--
-- Create Date:    
-- Design Name:    
-- Module Name:    k_2pi_sub - alg
-- Project Name:   
-- Target Device:  
-- Tool versions:  7.1i
--
-- === Brief description ===
--
-- M�dulo que resta a la entrada el valor 2*pi, aunque el formato del pipeline tenga una magnitud
-- limitada que no permita representar la constante 2*pi.
--
-- === Description ===
--
-- El uso habitual de esta entidad es en aquellos casos en los que se quiere mantener 0 <= |phi| <
-- PI, mediante la resta de la constante 2*pi en cuanto se detecte que el �ngulo phi acabe de
-- superar el l�mite superior de pi, pero se dispone de un pipeline con magnitud limitada. Con un
-- elemento restador del ancho del pipeline y una constante en una de sus entradas, no ser�a posible
-- realizar la resta.
--
-- Este bloque se encarga de internamente extender el pipeline, si es necesario, para representar la
-- constante 2*pi, y llevar a cabo la resta. 
--
-- == Necesidad ==
--
-- La codificaci�n elegida originalmente (FX3.16) obligaba a la utilizaci�n de este elemento, ya que
-- 2*pi no era un valor representable en el pipeline. Para comodidad, en lugar de "anchear" el
-- pipeline temporalmente en el punto donde fuese necesario el reajuste del valor de determinado
-- �ngulo, se dise�o este bloque.
--
-- Ahora mismo, el ancho de pipeline es 100% flexible. Las primeras pruebas nos parecen indicar que
-- al menos deberemos usar un FX4.16 o incluso FX5.16 (con tan s�lo 9 bits para la parte
-- fraccionaria), todas con capacidad para representar 2*pi. Este bloque parecer�a carecer de uso
--
-- Preferimos sin embargo mantener la t�ctica de que todos los �ngulos vayan en argumento principal
-- (-180 < 0 <= 180), y seguimos utilizando este elemento.
-- 
-- === TODO ===
--
-- == Check if constant adder is using "simplified logic" ==
--
-- 1.- A 17 bit adder is CORRECTLY inferred. But I'M ADDING A CONSTANT.
--      Check in the final implementation is design is simplified with k in mind.
--
-- === Revision ===
--
-- Revision 0.02 - Reworked: adapted to new to_vector and to_integer system, and made it
-- automatically detect if pipeline width must be extended.
--
-- Revision 0.01 - File Created
--------------------------------------------------------------------------------
library IEEE;
use WORK.COMMON.all;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity k_2pi_sub is
	generic (
		width : natural := PIPELINE_WIDTH;
                prec : natural := PIPELINE_PREC);
	port (
		i : in std_logic_vector(width - 1 downto 0);
		en : in std_logic;
		o : out std_logic_vector(width - 1 downto 0));
end k_2pi_sub;

architecture beh of k_2pi_sub is
        constant magn_size : natural := PIPELINE_WIDTH - PIPELINE_PREC - 1;
begin
        extended_generate : if magn_size < min_magn_size(TWO_PI) generate
        begin
                sub : process(i, en)
                        variable big_in, big_res : std_logic_vector(min_magn_size(TWO_PI) + 1 + PIPELINE_PREC downto 0);
                begin
                        big_in(width - 1 downto 0) := i;
                        big_in(big_in'high downto width) := (others => i(width - 1)); -- Sign extension
                        big_res := std_logic_vector(signed(big_in) + signed(to_vector(MINUS_TWO_PI, big_res'length, PIPELINE_PREC)));
                        if (en = '1') then
                                o(width - 2 downto 0) <= big_res(width - 2 downto 0);
                                o(width - 1) <= big_res(width); -- SIGN
                                                                -- EXTENSION
                                                                -- (compression :)
                        else
                                o <= i;
                        end if;
                end process;
        end generate;

        normal_generate : if magn_size >= min_magn_size(TWO_PI) generate
        begin
                sub : process(i, en)
                begin
                        if (en = '1') then
                                o <= std_logic_vector(signed(i) + signed(to_vector(MINUS_TWO_PI, width, prec)));
                        else
                                o <= i;
                        end if;
                end process;
        end generate;
end beh;
